package datatypes;
import FixedPoint::*;

`define IMG 8

typedef FixedPoint#(20,12) DataType;
typedef FixedPoint#(8,32) CoeffType;
typedef UInt#(16) ImgWidth;

endpackage
